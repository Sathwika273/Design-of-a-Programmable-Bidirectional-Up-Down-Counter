// Code your testbench here
// or browse Examples
`include "base.sv"
`include "generator.sv"
`include "interface.sv"
`include "driver.sv"
`include "monitor1.sv"
`include "monitor2.sv"
`include "scoreboard.sv"
`include "environment.sv"
`include "test.sv"
`include "top.sv"
